[%! "mux-entity.intralisp" %]
[% mux:config "s-mux" (mux:entity) %]
