[%! "mux-tb.intralisp" %]
[% let ((mux:data-lines 4) (mux:select-lines 2))
   (mux:tb) %]
