[%! "b-logic-vector-tb.intralisp" %]
[% b-logic-vector:tb %]
