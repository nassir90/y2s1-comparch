[%! "register-tb.intralisp" %]
[% register:tb %]
