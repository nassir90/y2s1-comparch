[%! "mux-entity.intralisp" %]
[% let ((mux:data-lines 16)
        (mux:select-lines 4))
 (mux:entity) %]
