[%! "b-logic-bit-entity.intralisp" %]
[% b-logic-bit:entity %]
