[%! "s-mux-tb.intralisp" %]
[% s-mux:tb %]
