[%! "b-logic-bit-tb.intralisp" %]
[% b-logic-bit:tb %]
