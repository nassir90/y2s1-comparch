[%! "memory-tb.intralisp" %]
[% memory:tb %]
