[%! "full-adder-entity.intralisp" %]
[% full-adder:entity %]
