[%! "functional-unit-tb.intralisp" %]
[% functional-unit:tb %]
