[%! "register-file-tb.intralisp" %]
[% register-file:tb %]
