[%! "mux-entity.intralisp" %]
[% let ((mux:size 1) (mux:data-lines 3) (mux:select-lines 2))
 (mux:entity)%]
