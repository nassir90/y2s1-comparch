[%! "pc-tb.intralisp" %]
[% pc:tb %]
