[%! "mux-entity.intralisp" %]
[% mux:config "cpu-2-17" (mux:entity) %]
