[%! "processor-1-entity.intralisp" %]
[% processor-1:entity %]
