[%! "mux-entity.intralisp" %]
[% mux:config "cpu-2-32" (mux:entity) %]
