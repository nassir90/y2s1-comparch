[%! "mux-tb.intralisp" %]
[% mux:config "cpu-2-32" (mux:tb) %]
