[%! "mux-entity.intralisp" %]
[% let ((mux:data-lines 3)
        (mux:select-lines 2))
 (mux:entity) %]
