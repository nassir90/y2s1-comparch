[%! "pc-entity.intralisp" %]
[% pc:entity %]
