[%! "flip-flop-tb.intralisp" %]
[% flip-flop:tb %]
