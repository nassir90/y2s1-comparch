[%! "logic-bitslice-entity.intralisp" %]
[% logic-bitslice:entity %]
