[%! "shifter-entity.intralisp" %]
[% shifter:entity %]
