[%! "logic-bit-entity.intralisp" %]
[% logic-bit:entity %]
