[%! "processor-entity.intralisp" %]
[% in-package :processor %]
[% processor:entity %]
