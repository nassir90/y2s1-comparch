[%! "b-logic-tb.intralisp" %]
[% b-logic:tb %]
