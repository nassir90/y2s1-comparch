[%! "decoder-tb.intralisp" %]
[% let ((decoder:output-lines 16)
        (decoder:input-lines 4))
 (decoder:tb) %]
