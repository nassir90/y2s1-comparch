[%! "sign-extend-entity.intralisp" %]
[% sign-extend:entity %]
