[%! "ripple-carry-adder-tb.intralisp" %]
[% ripple-carry-adder:tb %]
