[%! "mux-entity.intralisp" %]
[% mux:config "dp-3-1" (mux:entity) %]
