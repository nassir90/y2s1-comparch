[%! "datapath-entity.intralisp" %]
[% datapath:entity %]
