[%! "processor-2-entity.intralisp" %]
[% processor-2:entity %]
