[%! "mux-entity.intralisp" %]
[% mux:config "shifter-cflag" (mux:entity) %]
