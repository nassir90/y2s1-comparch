[%! "memory-entity.intralisp" %]
[% memory:entity %]
