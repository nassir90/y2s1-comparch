[%! "register-entity.intralisp" %]
[% let ((register:size 32)) (register:entity) %]
