[%! "control-memory-tb.intralisp" %]
[% control-memory:tb %]
