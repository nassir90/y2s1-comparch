[%! "zero-fill-entity.intralisp" %]
[% zero-fill:entity %]
