[%! "logic-vector-tb.intralisp" %]
[% logic-vector:tb %]
