[%! "datapath-tb.intralisp" %]
[% datapath:tb %]
