[%! "register-file-entity.intralisp" %]
[% register-file:entity %]
