[%! "logic-bitslice-tb.intralisp" %]
[% logic-bitslice:tb %]
