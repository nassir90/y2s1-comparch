[%! "mux-tb.intralisp" %]
[% mux:config "shifter-cflag" (mux:tb) %]
