[%! "status-register-tb.intralisp" %]
[% status-register:tb %]
