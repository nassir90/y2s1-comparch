[%! "mux-entity.intralisp" %]
[% let ((mux:size 1) (mux:data-lines 2) (mux:select-lines 1))
 (mux:entity)%]
