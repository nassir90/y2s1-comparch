[%! "alu-tb.intralisp" %]
[% alu:tb %]
