[%! "test-register-file-entity.intralisp" %]
[% test-register-file:entity %]
