[%! "test-register-file-tb.intralisp" %]
[% test-register-file:tb %]
