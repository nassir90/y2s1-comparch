[%! "ir-entity.intralisp" %]
[% ir:entity %]
