[%! "decoder-entity.intralisp" %]
[% let ((decoder:output-lines 32)
        (decoder:input-lines 5))
 (decoder:entity) %]
