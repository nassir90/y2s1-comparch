[%! "ir-tb.intralisp" %]
[% ir:tb %]
