[%! "processor-3-entity.intralisp" %]
[% processor-3:entity %]
