[%! "mux-entity.intralisp" %]
[% let ((mux:data-lines 32)
        (select-lines 5))
 (mux:entity) %]
