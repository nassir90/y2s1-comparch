[%! "zero-fill-tb.intralisp" %]
[% zero-fill:tb %]
