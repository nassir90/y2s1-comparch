[%! "b-logic-vector-entity.intralisp" %]
[% b-logic-vector:entity %]
