[%! "logic-vector-entity.intralisp" %]
[% logic-vector:entity %]
