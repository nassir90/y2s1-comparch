[%! "mux-entity.intralisp" %]
[% let ((mux:data-lines 4) (mux:select-lines 2) (mux:size 1))
   (mux:entity) %]
