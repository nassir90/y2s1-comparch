[%! "functional-unit-entity.intralisp" %]
[% functional-unit:entity %]
