[%! "b-logic-entity.intralisp" %]
[% b-logic:entity %]
