[%! "sign-extend-tb.intralisp" %]
[% sign-extend:tb %]
