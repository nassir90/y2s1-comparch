[%! "zero-detector-entity.intralisp" %]
[% zero-detector:entity %]
