[%! "shifter-tb.intralisp" %]
[% shifter:tb %]

