[%! "logic-bit-tb.intralisp" %]
[% logic-bit:tb %]
