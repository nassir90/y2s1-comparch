[%! "flip-flop-entity.intralisp" %]
[% flip-flop:entity %]
