[%! "car-entity.intralisp" %]
[% in-package :car %]
[% car:entity %]
