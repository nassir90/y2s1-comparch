[%! "processor-tb.intralisp" %]
[% processor:tb %]
