[%! "processor-3-tb.intralisp" %]
[% processor-3:tb %]
