[%! "mux-tb.intralisp" %]
[% let ((mux:data-lines 32)
        (select-lines 5))
 (mux:tb) %]
