[%! "mux-tb.intralisp" %]
[% mux:config "s-mux" (mux:tb) %]
