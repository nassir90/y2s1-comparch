[%! "processor-4-tb.intralisp" %]
[% processor-4:tb %]
