[%! "processor-4-entity.intralisp" %]
[% processor-4:entity %]
