[%! "car-tb.intralisp" %]
[% in-package :car %]
[% car:tb %]
