[%! "mux-tb.intralisp" %]
[% mux:config "cpu-2-17" (mux:tb) %]
