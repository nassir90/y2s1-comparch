[%! "zero-detector-tb.intralisp" %]
[% zero-detector:tb %]
