[%! "status-register-entity.intralisp" %]
[% status-register:entity %]
