[%! "mux-entity.intralisp" %]
[% let ((mux:data-lines 2) (mux:select-lines 1))
   (mux:entity) %]
