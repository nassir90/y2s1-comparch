[%! "mux-entity.intralisp" %]
[% mux:config "dp-cflag" (mux:entity) %]
