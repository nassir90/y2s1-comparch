[%! "ripple-carry-adder-entity.intralisp" %]
[% ripple-carry-adder:entity %]
