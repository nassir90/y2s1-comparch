[%! "processor-2-tb.intralisp" %]
[% processor-2:tb %]
