[%! "mux-tb.intralisp" %]
[% mux:config "dp-3-1" (mux:tb) %]
