[%! "s-mux-entity.intralisp" %]
[% s-mux:entity %]
