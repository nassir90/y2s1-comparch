[%! "alu-entity.intralisp" %]
[% alu:entity %]
