[%! "full-adder-tb.intralisp" %]
[% full-adder:tb %]
