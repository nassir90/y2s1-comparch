[%! "mux-tb.intralisp" %]
[% mux:config "dp-cflag" (mux:tb) %]
