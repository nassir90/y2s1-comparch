[%! "processor-1-tb.intralisp" %]
[% processor-1:tb %]
