[%! "control-memory-entity.intralisp" %]
[% control-memory:entity %]
